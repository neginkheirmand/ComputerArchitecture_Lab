library ieee; 
use ieee.std_logic_1164.all;
 entity fullAdder_tb is end entity fullAdder_tb; 
architecture test of fullAdder_tb is component full_adder is Port( i0, i1, cin: in std_logic; s, cout : out std_logic ); 
end component; 
signal in0   :std_logic;
signal in1   :std_logic; 
signal cin1  :std_logic; 
signal s1    :std_logic; 
signal cout1 :std_logic; 
begin FA:full_adder port map ( i0 => in0,  i1 => in1, cin => cin1, s => s1, cout => cout1); 
in0 <= '0', '1' after 100 ns, '0' after 200 ns; 
in1 <= '0', '0' after 100 ns, '1' after 200 ns; 
cin1 <= '0', '1' after 100 ns, '1' after 200 ns; 
end test;